module SCORE_DATA(clk_25MHz,count,data,data_adrs,score_t);
input clk_25MHz;
input [4:0] data_adrs;
input [3:0] count;
output reg [0:19] data;
output reg [0:99] score_t;
always @(posedge clk_25MHz)
begin
    case(count)
    4'd0:
        begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000011000000000;
        5'd03:data<=20'b00000011111111000000;
        5'd04:data<=20'b00000111111111100000;
        5'd05:data<=20'b00001111111111110000;
        5'd06:data<=20'b00001111111111110000;
        5'd07:data<=20'b00011111000011111000;
        5'd08:data<=20'b00011110000011111000;
        5'd09:data<=20'b00011110000001111000;
        5'd10:data<=20'b00111110000001111000;
        5'd11:data<=20'b00111110000001111000;
        5'd12:data<=20'b00111110000001111100;
        5'd13:data<=20'b00111100000001111100;
        5'd14:data<=20'b00111100000001111100;
        5'd15:data<=20'b00111100000001111100;
        5'd16:data<=20'b00111100000001111100;
        5'd17:data<=20'b00111100000001111100;
        5'd18:data<=20'b00111100000001111100;
        5'd19:data<=20'b00111110000001111100;
        5'd20:data<=20'b00111110000001111000;
        5'd21:data<=20'b00111110000001111000;
        5'd22:data<=20'b00111110000001111000;
        5'd23:data<=20'b00111110000011111000;
        5'd24:data<=20'b00011111000011111000;
        5'd25:data<=20'b00011111100111110000;
        5'd26:data<=20'b00011111111111110000;
        5'd27:data<=20'b00001111111111100000;
        5'd28:data<=20'b00000111111111000000;
        5'd29:data<=20'b00000011111110000000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;    
        endcase
        end
    4'd1:begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000000000000000;
        5'd04:data<=20'b00000001111000000000;
        5'd05:data<=20'b00000011111000000000;
        5'd06:data<=20'b00000111111000000000;
        5'd07:data<=20'b00011111111000000000;
        5'd08:data<=20'b00011111111000000000;
        5'd09:data<=20'b00011101111000000000;
        5'd10:data<=20'b00011001111000000000;
        5'd11:data<=20'b00000001111000000000;
        5'd12:data<=20'b00000001111000000000;
        5'd13:data<=20'b00000001111000000000;
        5'd14:data<=20'b00000001111000000000;
        5'd15:data<=20'b00000001111000000000;
        5'd16:data<=20'b00000001111000000000;
        5'd17:data<=20'b00000001111000000000;
        5'd18:data<=20'b00000001111000000000;
        5'd19:data<=20'b00000001111000000000;
        5'd20:data<=20'b00000001111000000000;
        5'd21:data<=20'b00000001111000000000;
        5'd22:data<=20'b00000001111000000000;
        5'd23:data<=20'b00000001111000000000;
        5'd24:data<=20'b00000001111000000000;
        5'd25:data<=20'b00000001111100000000;
        5'd26:data<=20'b00011111111111100000;
        5'd27:data<=20'b00011111111111100000;
        5'd28:data<=20'b00011111111111100000;
        5'd29:data<=20'b00011111111111100000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
        end
    4'd2:
        begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000001111100000000;
        5'd03:data<=20'b00000111111111000000;
        5'd04:data<=20'b00011111111111100000;
        5'd05:data<=20'b00011111111111100000;
        5'd06:data<=20'b00011111111111110000;
        5'd07:data<=20'b00011100011111110000;
        5'd08:data<=20'b00011000001111110000;
        5'd09:data<=20'b00000000000111110000;
        5'd10:data<=20'b00000000000111110000;
        5'd11:data<=20'b00000000000111110000;
        5'd12:data<=20'b00000000000111110000;
        5'd13:data<=20'b00000000001111110000;
        5'd14:data<=20'b00000000001111100000;
        5'd15:data<=20'b00000000001111100000;
        5'd16:data<=20'b00000000011111000000;
        5'd17:data<=20'b00000000111111000000;
        5'd18:data<=20'b00000000111110000000;
        5'd19:data<=20'b00000001111100000000;
        5'd20:data<=20'b00000011111000000000;
        5'd21:data<=20'b00000111111000000000;
        5'd22:data<=20'b00001111110000000000;
        5'd23:data<=20'b00001111100000000000;
        5'd24:data<=20'b00011111000000000000;
        5'd25:data<=20'b00011111111111111000;
        5'd26:data<=20'b00111111111111111000;
        5'd27:data<=20'b00111111111111111000;
        5'd28:data<=20'b00011111111111111000;
        5'd29:data<=20'b00011111111111110000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
        end
    4'd3:
        begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000011000000000;
            5'd03:data<=20'b00000111111111000000;
            5'd04:data<=20'b00001111111111100000;
            5'd05:data<=20'b00011111111111100000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011100001111110000;
            5'd08:data<=20'b00010000000111110000;
            5'd09:data<=20'b00000000000111110000;
            5'd10:data<=20'b00000000000111110000;
            5'd11:data<=20'b00000000000111110000;
            5'd12:data<=20'b00000000000111110000;
            5'd13:data<=20'b00000000001111100000;
            5'd14:data<=20'b00000111111111000000;
            5'd15:data<=20'b00001111111110000000;
            5'd16:data<=20'b00001111111111000000;
            5'd17:data<=20'b00000111111111110000;
            5'd18:data<=20'b00000000011111110000;
            5'd19:data<=20'b00000000000111111000;
            5'd20:data<=20'b00000000000011111000;
            5'd21:data<=20'b00000000000011111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011111000;
            5'd24:data<=20'b00010000000111111000;
            5'd25:data<=20'b00111100001111111000;
            5'd26:data<=20'b00111111111111110000;
            5'd27:data<=20'b00111111111111100000;
            5'd28:data<=20'b00011111111111000000;
            5'd29:data<=20'b00001111111110000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
            endcase
        end
    4'd4:
    begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000011111100000;
        5'd04:data<=20'b00000000011111100000;
        5'd05:data<=20'b00000000111111100000;
        5'd06:data<=20'b00000000111111100000;
        5'd07:data<=20'b00000001111111100000;
        5'd08:data<=20'b00000001111111100000;
        5'd09:data<=20'b00000011110111100000;
        5'd10:data<=20'b00000011110111100000;
        5'd11:data<=20'b00000111100111100000;
        5'd12:data<=20'b00000111100111100000;
        5'd13:data<=20'b00001111000111100000;
        5'd14:data<=20'b00001111000111100000;
        5'd15:data<=20'b00011110000111100000;
        5'd16:data<=20'b00011110000111100000;
        5'd17:data<=20'b00111100000111100000;
        5'd18:data<=20'b00111100000111100000;
        5'd19:data<=20'b00111000000111100000;
        5'd20:data<=20'b00111111111111111100;
        5'd21:data<=20'b00111111111111111100;
        5'd22:data<=20'b00111111111111111100;
        5'd23:data<=20'b00111111111111111100;
        5'd24:data<=20'b00000000000111110000;
        5'd25:data<=20'b00000000000111100000;
        5'd26:data<=20'b00000000000111100000;
        5'd27:data<=20'b00000000000111100000;
        5'd28:data<=20'b00000000000111100000;
        5'd29:data<=20'b00000000000111100000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd5:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00001111111111100000;
            5'd04:data<=20'b00011111111111110000;
            5'd05:data<=20'b00011111111111110000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011111111111100000;
            5'd08:data<=20'b00011110000000000000;
            5'd09:data<=20'b00011110000000000000;
            5'd10:data<=20'b00011110000000000000;
            5'd11:data<=20'b00011110000000000000;
            5'd12:data<=20'b00011110000000000000;
            5'd13:data<=20'b00011111111100000000;
            5'd14:data<=20'b00011111111111000000;
            5'd15:data<=20'b00011111111111100000;
            5'd16:data<=20'b00011111111111110000;
            5'd17:data<=20'b00001100011111111000;
            5'd18:data<=20'b00000000000111111000;
            5'd19:data<=20'b00000000000011111000;
            5'd20:data<=20'b00000000000011111000;
            5'd21:data<=20'b00000000000011111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011111000;
            5'd24:data<=20'b00000000000111111000;
            5'd25:data<=20'b00011000001111110000;
            5'd26:data<=20'b00011111111111110000;
            5'd27:data<=20'b00011111111111100000;
            5'd28:data<=20'b00011111111111000000;
            5'd29:data<=20'b00001111111100000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd6:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00000000111111110000;
            5'd04:data<=20'b00000011111111110000;
            5'd05:data<=20'b00000011111111110000;
            5'd06:data<=20'b00000111111111110000;
            5'd07:data<=20'b00001111100000000000;
            5'd08:data<=20'b00001111000000000000;
            5'd09:data<=20'b00011111000000000000;
            5'd10:data<=20'b00011110000000000000;
            5'd11:data<=20'b00011110000000000000;
            5'd12:data<=20'b00011110000000000000;
            5'd13:data<=20'b00011110011111000000;
            5'd14:data<=20'b00011111111111110000;
            5'd15:data<=20'b00011111111111111000;
            5'd16:data<=20'b00111111111111111000;
            5'd17:data<=20'b00111111000011111100;
            5'd18:data<=20'b00111110000001111100;
            5'd19:data<=20'b00011110000001111100;
            5'd20:data<=20'b00011110000001111100;
            5'd21:data<=20'b00011110000001111100;
            5'd22:data<=20'b00011110000001111100;
            5'd23:data<=20'b00011110000001111100;
            5'd24:data<=20'b00011111000001111000;
            5'd25:data<=20'b00011111100011111000;
            5'd26:data<=20'b00001111111111111000;
            5'd27:data<=20'b00001111111111110000;
            5'd28:data<=20'b00000111111111100000;
            5'd29:data<=20'b00000001111110000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd7:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000000000000000;
            5'd03:data<=20'b00011111111111111000;
            5'd04:data<=20'b00111111111111111000;
            5'd05:data<=20'b00111111111111111000;
            5'd06:data<=20'b00111111111111111000;
            5'd07:data<=20'b00011111111111111000;
            5'd08:data<=20'b00000000000011111000;
            5'd09:data<=20'b00000000000011111000;
            5'd10:data<=20'b00000000000111110000;
            5'd11:data<=20'b00000000000111110000;
            5'd12:data<=20'b00000000000111110000;
            5'd13:data<=20'b00000000001111100000;
            5'd14:data<=20'b00000000001111100000;
            5'd15:data<=20'b00000000001111000000;
            5'd16:data<=20'b00000000011111000000;
            5'd17:data<=20'b00000000011111000000;
            5'd18:data<=20'b00000000111110000000;
            5'd19:data<=20'b00000000111110000000;
            5'd20:data<=20'b00000000111110000000;
            5'd21:data<=20'b00000001111100000000;
            5'd22:data<=20'b00000001111100000000;
            5'd23:data<=20'b00000011111100000000;
            5'd24:data<=20'b00000011111000000000;
            5'd25:data<=20'b00000011111000000000;
            5'd26:data<=20'b00000111110000000000;
            5'd27:data<=20'b00000111110000000000;
            5'd28:data<=20'b00000111110000000000;
            5'd29:data<=20'b00000111100000000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd8:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000001000000000;
            5'd03:data<=20'b00000011111111000000;
            5'd04:data<=20'b00000111111111100000;
            5'd05:data<=20'b00001111111111110000;
            5'd06:data<=20'b00011111101111111000;
            5'd07:data<=20'b00011111000011111000;
            5'd08:data<=20'b00011110000001111000;
            5'd09:data<=20'b00011110000001111000;
            5'd10:data<=20'b00011110000001111000;
            5'd11:data<=20'b00011111000011111000;
            5'd12:data<=20'b00011111000111110000;
            5'd13:data<=20'b00001111111111100000;
            5'd14:data<=20'b00001111111111100000;
            5'd15:data<=20'b00000111111111000000;
            5'd16:data<=20'b00000011111111000000;
            5'd17:data<=20'b00000111111111110000;
            5'd18:data<=20'b00001111101111110000;
            5'd19:data<=20'b00011111000111111000;
            5'd20:data<=20'b00011110000011111000;
            5'd21:data<=20'b00111110000001111100;
            5'd22:data<=20'b00111100000001111100;
            5'd23:data<=20'b00111100000001111100;
            5'd24:data<=20'b00111110000001111000;
            5'd25:data<=20'b00111111000011111000;
            5'd26:data<=20'b00011111111111111000;
            5'd27:data<=20'b00011111111111110000;
            5'd28:data<=20'b00001111111111100000;
            5'd29:data<=20'b00000011111111000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd9:
    begin
        case(data_adrs)
            5'd00:data<=20'b00000000000000000000;
            5'd01:data<=20'b00000000000000000000;
            5'd02:data<=20'b00000000011000000000;
            5'd03:data<=20'b00000011111111000000;
            5'd04:data<=20'b00000111111111100000;
            5'd05:data<=20'b00001111111111110000;
            5'd06:data<=20'b00011111111111110000;
            5'd07:data<=20'b00011111000011111000;
            5'd08:data<=20'b00111110000011111000;
            5'd09:data<=20'b00111110000001111000;
            5'd10:data<=20'b00111100000001111000;
            5'd11:data<=20'b00111100000001111000;
            5'd12:data<=20'b00111110000001111000;
            5'd13:data<=20'b00111110000001111000;
            5'd14:data<=20'b00111110000001111000;
            5'd15:data<=20'b00011111000111111000;
            5'd16:data<=20'b00011111111111111000;
            5'd17:data<=20'b00011111111111111000;
            5'd18:data<=20'b00001111111111111000;
            5'd19:data<=20'b00000011111001111000;
            5'd20:data<=20'b00000000000001111000;
            5'd21:data<=20'b00000000000001111000;
            5'd22:data<=20'b00000000000011111000;
            5'd23:data<=20'b00000000000011110000;
            5'd24:data<=20'b00000000000111110000;
            5'd25:data<=20'b00011000001111100000;
            5'd26:data<=20'b00011111111111100000;
            5'd27:data<=20'b00011111111111000000;
            5'd28:data<=20'b00011111111110000000;
            5'd29:data<=20'b00001111111000000000;
            5'd30:data<=20'b00000000000000000000;
            5'd31:data<=20'b00000000000000000000;
        endcase
    end
    4'd10:
    begin
        case(data_adrs)
        5'd00:data<=20'b00000000000000000000;
        5'd01:data<=20'b00000000000000000000;
        5'd02:data<=20'b00000000000000000000;
        5'd03:data<=20'b00000000000000000000;
        5'd04:data<=20'b00000000000000000000;
        5'd05:data<=20'b00000000000000000000;
        5'd06:data<=20'b00000000000000000000;
        5'd07:data<=20'b00000000000000000000;
        5'd08:data<=20'b00000000000000000000;
        5'd09:data<=20'b00000000000000000000;
        5'd10:data<=20'b00000000011111000000;
        5'd11:data<=20'b00000000011111000000;
        5'd12:data<=20'b00000000011111000000;
        5'd13:data<=20'b00000000011111000000;
        5'd14:data<=20'b00000000000000000000;
        5'd15:data<=20'b00000000000000000000;
        5'd16:data<=20'b00000000000000000000;
        5'd17:data<=20'b00000000000000000000;
        5'd18:data<=20'b00000000000000000000;
        5'd19:data<=20'b00000000000000000000;
        5'd20:data<=20'b00000000000000000000;
        5'd21:data<=20'b00000000000000000000;
        5'd22:data<=20'b00000000000000000000;
        5'd23:data<=20'b00000000011111000000;
        5'd24:data<=20'b00000000011111000000;
        5'd25:data<=20'b00000000011111000000;
        5'd26:data<=20'b00000000011111000000;
        5'd27:data<=20'b00000000000000000000;
        5'd28:data<=20'b00000000000000000000;
        5'd29:data<=20'b00000000000000000000;
        5'd30:data<=20'b00000000000000000000;
        5'd31:data<=20'b00000000000000000000;
        endcase
    end
    default:
        data<=0;    
    endcase
end
always @(posedge clk_25MHz)
begin
    case(data_adrs)
        5'd00:score_t<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        5'd01:score_t<=100'b0000000110000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000;
        5'd02:score_t<=100'b0000111111110000000000011111110000000000011111111100000000001111111110000000001111111111110000000000;
        5'd03:score_t<=100'b0001111111111000000001111111111100000000111111111110000000001111111111100000001111111111110000000000;
        5'd04:score_t<=100'b0011111111111000000011111111111110000001111111111111000000001111111111110000001111111111110000000000;
        5'd05:score_t<=100'b0011100000011000000011110000011110000011110000001111100000001110000011110000001111000000000000000000;
        5'd06:score_t<=100'b0111100000000000000111100000000110000111100000000011100000001110000001111000001110000000000000000000;
        5'd07:score_t<=100'b0111000000000000000111000000000000000111000000000011110000001110000001111000001110000000000000000000;
        5'd08:score_t<=100'b0111000000000000001111000000000000000111000000000001110000001110000000111000001110000000000000000000;
        5'd09:score_t<=100'b0111000000000000001110000000000000001111000000000001110000001110000000111000001110000000000000000000;
        5'd10:score_t<=100'b0111100000000000001110000000000000001110000000000001111000001110000000111000001110000000000000001100;
        5'd11:score_t<=100'b0111100000000000011110000000000000001110000000000000111000001110000000111000001110000000000000001110;
        5'd12:score_t<=100'b0011110000000000011100000000000000001110000000000000111000001110000001111000001110000000000000001110;
        5'd13:score_t<=100'b0011111000000000011100000000000000001110000000000000111000001110000001110000001110000000000000001110;
        5'd14:score_t<=100'b0001111110000000011100000000000000001110000000000000111000001110000111100000001111111111100000001110;
        5'd15:score_t<=100'b0000111111000000011100000000000000001110000000000000111000001111111111100000001111111111100000000000;
        5'd16:score_t<=100'b0000011111110000011100000000000000011110000000000000111000001111111110000000001111111111100000000000;
        5'd17:score_t<=100'b0000000111111000011100000000000000001110000000000000111000001111111111000000001111000000000000000000;
        5'd18:score_t<=100'b0000000011111000011100000000000000001110000000000000111000001110000111000000001110000000000000000000;
        5'd19:score_t<=100'b0000000000111100011100000000000000001110000000000000111000001110000011100000001110000000000000000000;
        5'd20:score_t<=100'b0000000000111100011100000000000000001110000000000000111000001110000011100000001110000000000000000000;
        5'd21:score_t<=100'b0000000000011100011110000000000000001110000000000001111000001110000001110000001110000000000000000000;
        5'd22:score_t<=100'b0000000000011100001110000000000000001110000000000001110000001110000001110000001110000000000000000000;
        5'd23:score_t<=100'b0000000000011100001110000000000000001111000000000001110000001110000001110000001110000000000000000000;
        5'd24:score_t<=100'b0000000000011100001111000000000000000111000000000011110000001110000001111000001110000000000000000000;
        5'd25:score_t<=100'b0000000000011100000111000000000010000111100000000011100000001110000000111000001110000000000000000000;
        5'd26:score_t<=100'b0110000000111000000111100000001110000111100000000111100000001110000000111000001110000000000000001110;
        5'd27:score_t<=100'b0111100001111000000011111000111110000011111000011111000000001110000000111100001111000000000000001110;
        5'd28:score_t<=100'b0111111111110000000011111111111100000001111111111110000000001110000000011100001111111111111000001110;
        5'd29:score_t<=100'b0011111111100000000001111111111000000000111111111100000000001110000000011100001111111111111000001110;
        5'd30:score_t<=100'b0001111111000000000000011111100000000000001111111000000000001110000000011100000111111111111000001110;
        5'd31:score_t<=100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    endcase
end
endmodule